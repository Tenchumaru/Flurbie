parameter NR= 4;

typedef logic[4:0] regind_t;
typedef integer unsigned regval_t;
typedef regval_t regfile_t[NR];

parameter regfile_t ZeroRegFile= '{NR{0}};
parameter Flags= NR - 1;
parameter PC= Flags - 1;

function regfile_t subst_in(input regval_t pc, input regfile_t registers);
	return '{0, registers[1], pc, registers[Flags]};
endfunction

// shift operation
parameter logic[1:0] None= 0;
parameter logic[1:0] Left= 1;
parameter logic[1:0] LogicalRight= 2;
parameter logic[1:0] ArithmeticRight= 3;
parameter logic[2:0] Add= 3'b100;

parameter regval_t Nop= 32'h80000000;

interface i_fetch_to_decode();

logic hold, is_pc_changing;
regval_t instruction;

modport fetch_out(
	input hold, is_pc_changing,
	output instruction
);

modport decode_in(
	input instruction,
	output hold, is_pc_changing
);

endinterface

interface i_decode_to_read();

regval_t pc, adjustment;
regind_t destination, left_register, right_register;
logic[3:0] operation;
logic[2:0] adjustment_operation;
logic hold, destination_is_memory, right_is_memory, has_flushed, is_valid;

modport decode_out(
	input hold,
	output pc, adjustment,
	output destination, left_register, right_register,
	output operation,
	output adjustment_operation,
	output destination_is_memory, right_is_memory, has_flushed, is_valid
);

modport read_in(
	input pc, adjustment,
	input destination, left_register, right_register,
	input operation,
	input adjustment_operation,
	input destination_is_memory, right_is_memory, has_flushed, is_valid,
	output hold
);

endinterface

interface i_read_to_execute();

regval_t pc, adjustment, left_value, right_value;
regind_t destination;
logic[3:0] operation;
logic[2:0] adjustment_operation;
logic hold, destination_is_memory, has_flushed, is_valid;

modport read_out(
	input hold,
	output pc, adjustment, left_value, right_value,
	output destination,
	output operation,
	output adjustment_operation,
	output destination_is_memory, has_flushed, is_valid
);

modport execute_in(
	input pc, adjustment, left_value, right_value,
	input destination,
	input operation,
	input adjustment_operation,
	input destination_is_memory, has_flushed, is_valid,
	output hold
);

endinterface

interface i_execute_to_write();

regval_t pc, adjustment, destination_value;
regind_t destination;
logic[3:0] flags;
logic hold, destination_is_memory, has_flushed, is_valid;

modport execute_out(
	input hold,
	output pc, adjustment, destination_value,
	output destination,
	output flags,
	output destination_is_memory, has_flushed, is_valid
);
modport write_in(
	input pc, adjustment, destination_value,
	input destination,
	input flags,
	input destination_is_memory, has_flushed, is_valid,
	output hold
);

endinterface
